module  VGA_Controller(
  //  Host Side
  iRed,
  iGreen,
  iBlue,
  oRequest,
  //  VGA Side
  oVGA_R,
  oVGA_G,
  oVGA_B,
  oVGA_H_SYNC,
  oVGA_V_SYNC,
  oVGA_SYNC,
  oVGA_BLANK,
  oVGA_CLOCK,
  H_Cont,
  V_Cont,
  //  Control Signal
  iCLK,
  iRST_N
);

`include "VGA_Param.h"

//  Host Side
input [9:0] iRed;
input [9:0] iGreen;
input [9:0] iBlue;
output  reg oRequest;
//  VGA Side
output  [9:0] oVGA_R;
output  [9:0] oVGA_G;
output  [9:0] oVGA_B;
output  reg oVGA_H_SYNC;
output  reg oVGA_V_SYNC;
output      oVGA_SYNC;
output      oVGA_BLANK;
output      oVGA_CLOCK;
output     [9:0] H_Cont;
output     [9:0] V_Cont;
//  Control Signal
input       iCLK;
input       iRST_N;

//  Internal Registers and Wires
reg [9:0] H_Cont;
reg [9:0] V_Cont;
reg [9:0] Cur_Color_R;
reg [9:0] Cur_Color_G;
reg [9:0] Cur_Color_B;
wire			mCursor_EN;
wire				mRed_EN;
wire				mGreen_EN;
wire				mBlue_EN;

assign	oVGA_BLANK	=	oVGA_H_SYNC & oVGA_V_SYNC;
assign	oVGA_SYNC	=	1'b0;
assign	oVGA_CLOCK	=	iCLK;

assign	oVGA_R	=	(	H_Cont>=X_START 	&& H_Cont<X_START+H_SYNC_ACT &&
						V_Cont>=Y_START 	&& V_Cont<Y_START+V_SYNC_ACT )
						?	iRed	:	0;
assign	oVGA_G	=	(	H_Cont>=X_START 	&& H_Cont<X_START+H_SYNC_ACT &&
						V_Cont>=Y_START 	&& V_Cont<Y_START+V_SYNC_ACT )
						?	iGreen	:	0;
assign	oVGA_B	=	(	H_Cont>=X_START 	&& H_Cont<X_START+H_SYNC_ACT &&
						V_Cont>=Y_START 	&& V_Cont<Y_START+V_SYNC_ACT )
						?	iBlue	:	0;



//	Pixel LUT Address Generator
always@(posedge iCLK or negedge iRST_N)
begin
	if(!iRST_N)
	oRequest	<=	0;
	else
	begin
		if(	H_Cont>=X_START-2 && H_Cont<X_START+H_SYNC_ACT-2 &&
			V_Cont>=Y_START && V_Cont<Y_START+V_SYNC_ACT )
		oRequest	<=	1;
		else
		oRequest	<=	0;
	end
end

//	H_Sync Generator, Ref. 25.175 MHz Clock
always@(posedge iCLK or negedge iRST_N)
begin
	if(!iRST_N)
	begin
		H_Cont		<=	0;
		oVGA_H_SYNC	<=	0;
	end
	else
	begin
		//	H_Sync Counter
		if( H_Cont < H_SYNC_TOTAL )
		H_Cont	<=	H_Cont+1;
		else
		H_Cont	<=	0;
		//	H_Sync Generator
		if( H_Cont < H_SYNC_CYC )
		oVGA_H_SYNC	<=	0;
		else
		oVGA_H_SYNC	<=	1;
	end
end

//	V_Sync Generator, Ref. H_Sync
always@(posedge iCLK or negedge iRST_N)
begin
	if(!iRST_N)
	begin
		V_Cont		<=	0;
		oVGA_V_SYNC	<=	0;
	end
	else
	begin
		//	When H_Sync Re-start
		if(H_Cont==0)
		begin
			//	V_Sync Counter
			if( V_Cont < V_SYNC_TOTAL )
			V_Cont	<=	V_Cont+1;
			else
			V_Cont	<=	0;
			//	V_Sync Generator
			if(	V_Cont < V_SYNC_CYC )
			oVGA_V_SYNC	<=	0;
			else
			oVGA_V_SYNC	<=	1;
		end
	end
end

endmodule